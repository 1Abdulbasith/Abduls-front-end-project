<svg xmlns="http://www.w3.org/2000/svg" width="564.8103" height="449.94076" viewBox="0 0 564.8103 449.94076" xmlns:xlink="http://www.w3.org/1999/xlink"><g><g><polygon points="496.1376 436.61569 484.39597 436.61456 478.81042 391.32495 496.13998 391.32614 496.1376 436.61569" fill="#ffb6b6"/><path d="M496.5509,448.86453l-36.10718-.00137v-.45657c.00052-7.76151,6.29242-14.05328,14.05392-14.05371h.00089l6.59543-5.0036,12.3056,5.00439,3.15192,.00006-.00058,14.5108Z" fill="#2f2e41"/></g><g><polygon points="444.08279 436.61569 432.34119 436.61456 426.75562 391.32495 444.08521 391.32614 444.08279 436.61569" fill="#ffb6b6"/><path d="M444.49609,448.86453l-36.10718-.00137v-.45657c.00052-7.76151,6.29242-14.05328,14.05392-14.05371h.00089l6.59543-5.0036,12.3056,5.00439,3.15192,.00006-.00058,14.5108Z" fill="#2f2e41"/></g><path d="M438.48767,183.86459l67.74255,1.42616s12.17853,19.96622,2.8804,48.13286l1.04156,7.84387-4.27847,12.12234-2.13925,37.08014,2.13925,5.70462-1.42615,10.6962s5.70462,70.59485-8.55695,106.24881l-17.11389-.71307-6.41772-93.02316,3.5654-6.80795-.71307-2.85233-8.55695-42.78476-8.55695,22.10547v12.28238l-7.84387,9.11002s2.85233,84.14334-4.99155,101.25726h-19.16049l-7.22345-114.09268,7.1308-66.31638-1.42615-4.27847,2.13925-2.13924-1.42615-7.13078,13.19196-33.87128-.00012-.00003Z" fill="#2f2e41"/><path d="M467.36737,53.72761l20.67929-4.99156,5.70462,13.54851s29.51471,15.68775,30.94092,37.08013c0,0,4,17.1139,.43457,24.95778-3.56543,7.84386-18.54007,32.80164-18.54007,32.80164,0,0,13.54849,43.49783,9.98312,45.63708s-88.42184-2.13924-88.42184-6.41771,14.12234-49.20247,14.12234-49.20247l2.99155-77.01257,19.25314-7.13079,2.85233-9.27003,.00003-.00002Z" fill="#3f3d56"/><path d="M522.49719,229.26281c-4.32812-2.18115-6.06903-7.45773-3.88818-11.78589,.21954-.43568,.47803-.83762,.75598-1.21933l-11.50684-78.89287,15.93066,.50961,8.33337,76.86882c3.02032,2.56178,4.02191,6.93852,2.16089,10.63158-2.18085,4.32817-7.45752,6.06889-11.78595,3.88808h.00006Z" fill="#ffb6b6"/><path d="M371.33841,192.02793c-1.74237-4.52263,.51102-9.60155,5.03342-11.34416,.45523-.17542,.91669-.29967,1.379-.39581l44.45221-66.18528,11.46213,11.07548-45.44449,62.55444c.5177,3.92645-1.67923,7.84212-5.53818,9.32889-4.52243,1.74261-9.60132-.511-11.34409-5.03355Z" fill="#ffb6b6"/><path d="M493.46826,117.46573c-4.50104-15.46355,2.97473-31.24023,19.07983-31.16403,4.65497,.02203,8.27142,1.3728,9.27374,5.11178,3.50812,13.08646,5.42102,32.8406,5.42102,32.8406l4.16156,21.0321-2.52063,4.36699,5.25488,14.09471-2.54901,6.66808-.55109,34.05193-12.83545-.71307-14.14221-25.95921-5.40778-3.21553s4.34204-41.972-4.29492-54.05681l-.88998-3.05752h.00003Z" fill="#3f3d56"/><path d="M435.97525,79.40956c7.50537-14.24957,26.72006-17.6249,38.25119-6.38149,3.33292,3.24976,4.99576,6.73378,3.11914,10.11948-6.56818,11.84994-21.793,24.60873-21.793,24.60873l-18.74896,30.1414-4.84686,1.38994-6.01218,13.7887-12.88364,15.14767-17.06436,8.99919-9.98312-9.98311,2.11987-12.83292,25.69025-34.23032s18.4845-23.25715,20.66769-37.94979l1.48398-2.81748v-.00002Z" fill="#3f3d56"/><path d="M471.29678,49.55995c.47229,.05676,.94308,.09937,1.41153,.12074,1.45734,.07992,2.89713-.00317,4.28467-.23844,4.21613-.67573,8.04633-2.67263,11.0018-5.60105,3.12457-3.09,5.26291-7.2143,5.84094-11.90953,1.35419-11.08279-6.53763-21.17844-17.62042-22.53263-10.92374-1.34261-20.8815,6.29773-22.47101,17.12611-.02499,.16763-.05075,.3282-.0687,.49507-1.35342,11.08988,6.53058,21.1792,17.62119,22.53972v.00002Z" fill="#ffb6b6"/><path d="M449.18701,25.78329c2.87085,1.41972,7.5618-3.04364,9.3584-.47564,.29178-.55496,.61414-1.09167,.93253-1.59923,.28821-.45416,.70035-1.42364,1.17737-1.58967-.60361,1.45626-.47043,3.42853,.15594,5.1183,2.83197,1.05813,6.53894-1.28412,9.16-4.05461,4.11569-4.34412,10.83603,6.7955,9.24701,12.56046,2.02228-2.46946,6.41068-1.07667,7.89767,1.74692,1.48627,2.81653-1.02509,5.07323-1.56219,8.2149l4.05411-.51486c2.55783-2.49121,2.37894-6.68905,4.48535-9.57637,3.51816-4.83207,4.88135-9.76236,2.23651-14.74927-2.34604-4.40945-2.56531-10.11622-6.86929-12.6584,1.88055-.91942-4.80698,.51694-3.02066-2.47936,1.79419-2.99001-7.76917-3.35292-8.39297-1.75104-2.73279-3.27058-5.48917-5.42694-8.85068-2.80627-3.30151,2.57832-2.95984,5.28843-6.83731,5.04556-1.8194-.11273-1.6196,3.27962-2.70126,4.75862-1.07535,1.4711-5.25543,2.41549-5.45883,2.25806-1.1041-.86381-4.86032,6.48971-4.86032,6.48971,0,0-3.04572,4.6235-.15134,6.06219h-.00003Z" fill="#2f2e41"/></g><path d="M196.15526,154.13037c67.93102,0,123.00002,55.06897,123.00002,123s-55.069,123-123.00002,123-161.94494-67.3513-123-123,55.06898-123,123-123Z" fill="#f2f2f2"/><path d="M360.7818,159.98167c-1.10303,0-2,.89697-2,2v64c0,1.10303,.89697,2,2,2s2-.89697,2-2v-64c0-1.10303-.89697-2-2-2Z" fill="#3f3d56"/><path d="M24.7818,111.98166c-1.10303,0-2,.89697-2,2v15.99999c0,1.10303,.89697,2,2,2s2-.89697,2-2v-16c0-1.10303-.89697-2-2-1.99999Z" fill="#3f3d56"/><path d="M24.7818,159.98167c-1.10303,0-2,.89697-2,2v31c0,1.10303,.89697,2,2,2s2-.89697,2-2v-31c0-1.10303-.89697-2-2-2Z" fill="#3f3d56"/><path d="M24.7818,203.98167c-1.10303,0-2,.89697-2,2v31c0,1.10303,.89697,2,2,2s2-.89697,2-2v-31c0-1.10303-.89697-2-2-2Z" fill="#3f3d56"/><path d="M204.15526,48.98167c-1.10303,0-2,.89697-2,2v31c0,1.10303,.89697,2,2,2s2-.89697,2-2v-31c0-1.10303-.89697-2-2-2Z" fill="#3f3d56"/><g><path d="M510.55136,432.60781c2.06595,.12936,3.20767-2.43738,1.64468-3.93332l-.15552-.61819c.02045-.0495,.04108-.09897,.06177-.14838,2.08923-4.98181,9.16992-4.94742,11.24139,.04178,1.83856,4.42816,4.17944,8.86389,4.7558,13.54593,.25836,2.0668,.14215,4.17236-.31647,6.20047,4.30804-9.41058,6.57513-19.68661,6.57513-30.02078,0-2.59653-.14215-5.19302-.43274-7.78296-.23901-2.11853-.56842-4.22409-.99469-6.31033-2.30573-11.27719-7.29852-22.01825-14.50012-30.98962-3.46198-1.89249-6.34906-4.85065-8.09296-8.39651-.6265-1.2789-1.1174-2.65463-1.34991-4.05618,.39398,.05167,1.48557-5.94867,1.18842-6.3168,.54907-.83316,1.53177-1.24734,2.13147-2.06033,2.9823-4.0434,7.09119-3.3374,9.23621,2.15726,4.58221,2.31265,4.62659,6.14807,1.81494,9.83682-1.78876,2.34683-2.03455,5.52234-3.60406,8.03479,.1615,.2067,.32947,.40695,.49091,.61365,2.96106,3.79788,5.52209,7.88,7.68103,12.16858-.61017-4.7662,.29065-10.50821,1.82642-14.20959,1.74817-4.21732,5.0249-7.76917,7.91046-11.41501,3.466-4.37924,10.57336-2.46805,11.18402,3.08331,.00592,.05374,.01166,.10745,.01733,.16119-.42859,.24179-.84851,.49866-1.25867,.76993-2.33948,1.54724-1.53094,5.17386,1.24109,5.60175l.06274,.00967c-.15503,1.54367-.41986,3.07443-.80731,4.57938,3.70178,14.3158-4.2901,19.52991-15.70148,19.76413-.25189,.12915-.49738,.25833-.74927,.3811,1.15619,3.25525,2.07983,6.59448,2.7644,9.97891,.61359,2.99042,1.03992,6.01318,1.27887,9.04889,.29718,3.83005,.2713,7.6796-.0517,11.50323l.01941-.13562c.82025-4.21115,3.10669-8.14462,6.42657-10.87027,4.94562-4.06265,11.9328-5.55869,17.26825-8.82425,2.56836-1.57196,5.85944,.45944,5.41119,3.43707l-.02179,.14261c-.79443,.32288-1.56946,.69754-2.31873,1.11734-.42859,.24185-.84845,.49866-1.25867,.76993-2.33948,1.5473-1.53094,5.17392,1.24109,5.60181l.06281,.00964c.04523,.00647,.08398,.01294,.12909,.01944-1.36279,3.23581-3.26166,6.23923-5.63855,8.82922-2.31464,12.49713-12.25604,13.68283-22.8902,10.04355h-.00647c-1.1626,5.06378-2.86127,10.01126-5.04437,14.7262h-18.0202c-.06464-.20023-.12274-.40692-.18088-.60718,1.66641,.10342,3.34573,.0065,4.9863-.29703-1.33704-1.64059-2.67395-3.2941-4.01096-4.93463-.03229-.03229-.05817-.06461-.08398-.09689-.67816-.8396-1.36282-1.67282-2.04099-2.51245l-.00037-.00101c-.04245-2.57755,.26651-5.14661,.87875-7.63983l.00058-.00034-.00009-.00006Z" fill="#f2f2f2"/><path d="M0,448.75076c0,.66003,.53003,1.19,1.19006,1.19H563.48004c.65997,0,1.19-.52997,1.19-1.19,0-.65997-.53003-1.19-1.19-1.19H1.19006c-.66003,0-1.19006,.53003-1.19006,1.19Z" fill="#ccc"/></g><path d="M142.37598,268.83935H73.15526v-2h69.2207c6.01318,0,10.90527-4.89258,10.90527-10.90625v-46.80273h2v46.80273c0,7.11621-5.78906,12.90625-12.90527,12.90625h.00002Z" fill="#dc1246"/><rect x="117.01903" y="370.29443" width="157.43605" height="2" fill="#dc1246"/><g><path d="M374.34299,255.466h-84.0918c-4.53809,0-8.22998-3.69189-8.22998-8.22998v-83.06592c0-4.53809,3.69189-8.22998,8.22998-8.22998h84.0918c4.53809,0,8.22998,3.69189,8.22998,8.22998v83.06592c0,4.53809-3.69189,8.22998-8.22998,8.22998Z" fill="#e6e6e6"/><path d="M305.91171,158.39219c-11.84012,0-21.43842,9.5983-21.43842,21.43842v65.64299c0,4.16435,3.37589,7.54022,7.54022,7.54022h51.41989c20.26184,0,36.68732-16.42548,36.68732-36.68733v-50.39409c0-4.16435-3.37589-7.54022-7.54022-7.54022h-66.66879v.00002Z" fill="#fff"/><g><path d="M354.81924,182.53161h-45.22061c-.86273,0-1.5647-.702-1.5647-1.56471s.702-1.56439,1.5647-1.56439h45.22061c.86273,0,1.56439,.70166,1.56439,1.56439s-.70166,1.56471-1.56439,1.56471Z" fill="#e6e6e6"/><path d="M354.81924,215.89521h-45.22061c-.86273,0-1.5647-.702-1.5647-1.56471s.702-1.56439,1.5647-1.56439h45.22061c.86273,0,1.56439,.70166,1.56439,1.56439s-.70166,1.56471-1.56439,1.56471Z" fill="#e6e6e6"/><path d="M373.1824,199.22434h-81.9469c-.86273,0-1.5647-.702-1.5647-1.56471s.702-1.56439,1.5647-1.56439h81.9469c.86273,0,1.56439,.70166,1.56439,1.56439s-.70166,1.56471-1.56439,1.56471Z" fill="#e6e6e6"/></g><path d="M374.01913,229.46084h-29.60361c-.86273,0-1.5647-.702-1.5647-1.56471s.702-1.56439,1.5647-1.56439h29.60361c.86273,0,1.56439,.70166,1.56439,1.56439s-.70166,1.56471-1.56439,1.56471Z" fill="#e6e6e6"/></g><g><path d="M197.71127,420.97035h-66.77454c-3.60355,0-6.53516-2.93161-6.53516-6.53516v-65.95993c0-3.60355,2.93161-6.53516,6.53516-6.53516h66.77457c3.60355,0,6.53516,2.93161,6.53516,6.53516v65.95993c0,3.60355-2.93161,6.53516-6.53516,6.53516h-.00002Z" fill="#e6e6e6"/><path d="M143.37224,343.88719c-9.40184,0-17.02355,7.6217-17.02355,17.02356v52.12497c0,3.30679,2.68067,5.98746,5.98745,5.98746h40.83086c16.08928,0,29.13222-13.04294,29.13222-29.1322v-40.0163c0-3.30679-2.68066-5.98746-5.98746-5.98746h-52.93953l.00002-.00003Z" fill="#fff"/><g><path d="M182.20811,363.05549h-35.9082c-.68506,0-1.24249-.55743-1.24249-1.24249s.55742-1.24222,1.24249-1.24222h35.9082c.68506,0,1.24223,.55716,1.24223,1.24222s-.55717,1.24249-1.24223,1.24249Z" fill="#e6e6e6"/><path d="M182.20811,389.54847h-35.9082c-.68506,0-1.24249-.55743-1.24249-1.24249s.55742-1.24222,1.24249-1.24222h35.9082c.68506,0,1.24223,.55716,1.24223,1.24222s-.55717,1.24249-1.24223,1.24249Z" fill="#e6e6e6"/><path d="M196.78969,376.31068h-65.07135c-.68506,0-1.24249-.55743-1.24249-1.24249s.55742-1.24222,1.24249-1.24222h65.07135c.68506,0,1.24223,.55716,1.24223,1.24222s-.55717,1.24249-1.24223,1.24249Z" fill="#e6e6e6"/></g><path d="M197.4541,400.32048h-23.50725c-.68506,0-1.24249-.55743-1.24249-1.24249s.55742-1.24222,1.24249-1.24222h23.50725c.68506,0,1.24223,.55716,1.24223,1.24222s-.55717,1.24249-1.24223,1.24249Z" fill="#e6e6e6"/></g><g><path d="M151.04003,208.62567h-49.3827c-2.66499,0-4.83304-2.16805-4.83304-4.83303v-48.78026c0-2.66498,2.16805-4.83303,4.83303-4.83303h49.38271c2.66498,0,4.83303,2.16805,4.83303,4.83303v48.78026c0,2.66498-2.16805,4.83303-4.83303,4.83303h-.00001Z" fill="#e6e6e6"/><path d="M110.85394,151.6193c-6.95307,0-12.58966,5.63658-12.58966,12.58967v38.5487c0,2.44552,1.98247,4.42799,4.42798,4.42799h30.19621c11.89873,0,21.54455-9.64582,21.54455-21.54454v-29.5938c0-2.44552-1.98247-4.42799-4.42799-4.42799h-39.1511v-.00002Z" fill="#fff"/><g><path d="M139.57477,165.7951h-26.55569c-.50663,0-.91888-.41225-.91888-.91888s.41224-.91867,.91888-.91867h26.55569c.50663,0,.91869,.41204,.91869,.91867s-.41206,.91888-.91869,.91888Z" fill="#e6e6e6"/><path d="M139.57477,185.38782h-26.55569c-.50663,0-.91888-.41225-.91888-.91888s.41224-.91867,.91888-.91867h26.55569c.50663,0,.91869,.41204,.91869,.91867s-.41206,.91888-.91869,.91888Z" fill="#e6e6e6"/><path d="M150.35848,175.59789h-48.12311c-.50663,0-.91888-.41225-.91888-.91888s.41224-.91867,.91888-.91867h48.12311c.50663,0,.91869,.41204,.91869,.91867s-.41206,.91888-.91869,.91888Z" fill="#e6e6e6"/></g><path d="M150.84984,193.35418h-17.38464c-.50663,0-.91888-.41225-.91888-.91888s.41224-.91867,.91888-.91867h17.38464c.50663,0,.91869,.41204,.91869,.91867s-.41206,.91888-.91869,.91888Z" fill="#e6e6e6"/></g><circle cx="295.15527" cy="260.13037" r="10" fill="#dc1246"/><circle cx="154.15526" cy="209.13035" r="10" fill="#dc1246"/><circle cx="202.15526" cy="346.13037" r="10" fill="#dc1246"/><g><ellipse cx="223.75633" cy="66.65212" rx="12.46327" ry="12.20069" fill="#f2f2f2"/><path d="M323.66919,62.47819h-67.08496c-2.30142,0-4.17392-1.87249-4.17392-4.17392s1.8725-4.17392,4.17392-4.17392h67.08496c2.30142,0,4.17392,1.87249,4.17392,4.17392s-1.8725,4.17392-4.17392,4.17392Z" fill="#f2f2f2"/><path d="M376.02252,76.6053h-119.43829c-2.30142,0-4.17392-1.87249-4.17392-4.17392s1.8725-4.17392,4.17392-4.17392h119.43829c2.30142,0,4.17392,1.87249,4.17392,4.17392s-1.8725,4.17392-4.17392,4.17392Z" fill="#f2f2f2"/></g><g><ellipse cx="43.35911" cy="122.23425" rx="8.06605" ry="7.8961" fill="#f2f2f2"/><path d="M108.02125,119.53295h-43.4164c-1.48945,0-2.7013-1.21185-2.7013-2.7013s1.21185-2.7013,2.7013-2.7013h43.4164c1.48945,0,2.7013,1.21185,2.7013,2.7013s-1.21185,2.7013-2.70129,2.7013Z" fill="#f2f2f2"/><path d="M141.90355,128.67582H64.60485c-1.48945,0-2.7013-1.21185-2.7013-2.7013s1.21185-2.7013,2.7013-2.7013h77.2987c1.48946,0,2.70129,1.21185,2.70129,2.7013s-1.21185,2.7013-2.70129,2.7013Z" fill="#f2f2f2"/></g><g><ellipse cx="285.3591" cy="403.23425" rx="8.06604" ry="7.89609" fill="#f2f2f2"/><path d="M350.02124,400.53295h-43.41641c-1.48944,0-2.70129-1.21185-2.70129-2.70129s1.21185-2.70129,2.70129-2.70129h43.41641c1.48944,0,2.70129,1.21185,2.70129,2.70129s-1.21185,2.70129-2.70129,2.70129Z" fill="#f2f2f2"/><path d="M383.90356,409.67581h-77.29871c-1.48944,0-2.70129-1.21185-2.70129-2.70129s1.21185-2.70129,2.70129-2.70129h77.29871c1.48944,0,2.70129,1.21185,2.70129,2.70129s-1.21185,2.70129-2.70129,2.70129Z" fill="#f2f2f2"/></g><rect x="186.40511" y="155.97038" width="2" height="95" fill="#e6e6e6"/><circle cx="187.40511" cy="250.97038" r="6.00001" fill="#e6e6e6"/><circle cx="278.40511" cy="319.97039" r="6" fill="#e6e6e6"/><circle cx="116.40511" cy="237.97038" r="6" fill="#e6e6e6"/><rect x="81.39766" y="238.47578" width="32.82787" height="2.00092" transform="translate(-7.20166 3.0694) rotate(-1.73401)" fill="#e6e6e6"/><polygon points="327.21616 342.94012 277.4603 342.94012 277.4603 319.97039 279.4603 319.97039 279.4603 340.94012 327.21616 340.94012 327.21616 342.94012" fill="#e6e6e6"/><circle cx="113.94232" cy="303.48553" r="6" fill="#e6e6e6"/><polygon points="162.16098 326.45526 112.40511 326.45526 112.40511 303.48553 114.40511 303.48553 114.40511 324.45526 162.16098 324.45526 162.16098 326.45526" fill="#e6e6e6"/><rect x="75.42269" y="280.65496" width="238.98243" height="2" fill="#e6e6e6"/></svg>
